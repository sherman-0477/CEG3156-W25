library verilog;
use verilog.vl_types.all;
entity FPMult_vlg_vec_tst is
end FPMult_vlg_vec_tst;
